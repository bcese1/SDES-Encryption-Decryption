----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 
-- Design Name: 
-- Module Name: EP - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity EP is
    Port ( input : in STD_LOGIC_VECTOR (3 downto 0);
           expanded : out STD_LOGIC_VECTOR (7 downto 0));
end EP;

architecture Behavioral of EP is

begin

expanded(0) <= input(3);
expanded(1) <= input(0);
expanded(2) <= input(1);
expanded(3) <= input(2);
expanded(4) <= input(1);
expanded(5) <= input(2);
expanded(6) <= input(3);
expanded(7) <= input(0);

end Behavioral;
